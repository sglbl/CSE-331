library verilog;
use verilog.vl_types.all;
entity testbench_cypher_detect is
end testbench_cypher_detect;
