library verilog;
use verilog.vl_types.all;
entity testbench_control is
end testbench_control;
