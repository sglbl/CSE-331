module sll(input [15:0] a, input [15:0] b, input [3:0] shamt, output [15:0] result);

    wire [15:0] temp;
    wire [15:0] temp2;


endmodule